library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity programa_helloworld_int_FLIP is
	port( address : in std_logic_vector(7 downto 0);
		clk : in std_logic;
		dout : out std_logic_vector(15 downto 0));
	end;

architecture v1 of programa_helloworld_int_FLIP is

	constant ROM_WIDTH: INTEGER:= 16;
	constant ROM_LENGTH: INTEGER:= 256;

	subtype rom_word is std_logic_vector(ROM_WIDTH-1 downto 0);
	type rom_table is array (0 to ROM_LENGTH-1) of rom_word;

constant rom: rom_table := rom_table'(
	"1111000000000000",
	"1101100001100111",
	"0000000101001001",
	"1101100001110100",
	"0000000101101110",
	"1101100001110100",
	"0000000101110100",
	"1101100001110100",
	"0000000101110010",
	"1101100001110100",
	"0000000101101111",
	"1101100001110100",
	"0000000101100100",
	"1101100001110100",
	"0000000101110101",
	"1101100001110100",
	"0000000101111010",
	"1101100001110100",
	"0000000101100011",
	"1101100001110100",
	"0000000101100001",
	"1101100001110100",
	"0000000100100000",
	"1101100001110100",
	"0000000101110101",
	"1101100001110100",
	"0000000101101110",
	"1101100001110100",
	"0000000100100000",
	"1101100001110100",
	"0000000101100011",
	"1101100001110100",
	"0000000101100001",
	"1101100001110100",
	"0000000101110010",
	"1101100001110100",
	"0000000110100000",
	"1101100001110100",
	"0000000101100011",
	"1101100001110100",
	"0000000101110100",
	"1101100001110100",
	"0000000101100101",
	"1101100001110100",
	"0000000101110010",
	"1101100001110100",
	"0000000100111010",
	"1101100001110100",
	"0000000100100000",
	"1101100001110100",
	"1101100001100111",
	"0100011001000000",
	"0000000101111000",
	"1101100001110100",
	"0000000100111101",
	"1101100001110100",
	"0100000111000000",
	"1101100001110100",
	"0000000100100000",
	"1101100001110100",
	"0000000101000011",
	"1101100001110100",
	"0000000101001111",
	"1101100001110100",
	"0000000101001101",
	"1101100001110100",
	"0000000100110010",
	"1101100001110100",
	"0000000100101000",
	"1101100001110100",
	"0000000101111000",
	"1101100001110100",
	"0000000100101111",
	"1101100001110100",
	"0000000100110001",
	"1101100001110100",
	"0000000100110101",
	"1101100001110100",
	"0000000100101001",
	"1101100001110100",
	"0000000100111101",
	"1101100001110100",
	"1000111001000011",
	"1101100010001000",
	"1101100010001000",
	"1101100010001000",
	"1101100010001000",
	"1101100010001000",
	"1101100010001000",
	"1101100010001000",
	"1000011101000011",
	"0100011011100000",
	"1010111000000000",
	"0100000111000000",
	"1101100001110100",
	"0000000100001010",
	"1101100001110100",
	"1101000000000001",
	"0000011000001001",
	"0011011000000001",
	"1101010101100011",
	"0000011000001001",
	"1101000001100011",
	"1000001011111111",
	"0000101010000000",
	"1101010101100111",
	"1101100010001000",
	"0000001100001001",
	"1101100010000001",
	"1010001000001110",
	"1000000011111111",
	"0000100010000000",
	"0101001000000000",
	"0011001100000001",
	"1101010101101100",
	"1001000000000000",
	"0000000000000000",
	"1000100011111111",
	"1101100010000001",
	"0000001100001000",
	"1000100111111111",
	"1101100010000001",
	"1010000100001110",
	"0011001100000001",
	"1101010101111000",
	"0000000011111111",
	"1000100011111111",
	"1101100010000001",
	"1001000000000000",
	"0000010000000011",
	"0000010100100010",
	"0011010100000001",
	"1101010110000011",
	"0011010000000001",
	"1101010110000010",
	"1001000000000000",
	"0000010000000011",
	"0000010100010000",
	"0011010100000001",
	"1101010110001010",
	"0011010000000001",
	"1101010110001001",
	"1001000000000000",
	"1111000000000000",
	"1101100001100111",
	"1111101000000000",
	"0100000101000000",
	"1101100001110100",
	"0010011000110000",
	"0100000111000000",
	"1101100001110100",
	"1011000000000001",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"1101000010001111");

begin

process (clk)
begin
	if clk'event and clk = '1' then
		dout <= rom(conv_integer(address));
	end if;
end process;
end v1;
